module implicit(a,b,out);
  input a,b;
  assign out=a|b;
endmodule
