module multiple_initial;
  reg clk,a,b,c,e,d;
  initial clk=0; 
  initial a=0;
  initial b=0;
  initial c=0;
  initial d=0;
  initial d=0;
endmodule
